module boolean_function_1(
input A,
input B,
output F);

assign F= ~A & ~B;
endmodule